interface myBus;

        logic           a;
        logic           b;
        logic   [7:0]   c;

endinterface
